`ifndef RKV_AHBRAM_ELEMENT_SEQUENCES_SVH
`define RKV_AHBRAM_ELEMENT_SEQUENCES_SVH

`include "rkv_ahbram_base_element_sequence.sv"
`include "rkv_ahbram_single_read_seq.sv"
`include "rkv_ahbram_single_write_seq.sv"

`endif//RKV_AHBRAM_ELEMENT_SEQUENCES_SVH
