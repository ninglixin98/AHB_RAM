`ifndef LVC_AHB_PKG_SV
`define LVC_AHB_PKG_SV

package lvc_ahb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "lvc_ahb_defines.svh"
  `include "lvc_ahb_types.sv"
  `include "lvc_ahb_configuration.sv"
  `include "lvc_ahb_agent_configuration.sv"
  `include "lvc_ahb_transaction.sv" 
  `include "lvc_ahb_sequencer.sv"
  `include "lvc_ahb_driver.sv"
  `include "lvc_ahb_monitor.sv"
  `include "lvc_ahb_master_transaction.sv"
  `include "lvc_ahb_master_driver.sv"
  `include "lvc_ahb_master_monitor.sv"
  `include "lvc_ahb_master_sequencer.sv"
  `include "lvc_ahb_master_agent.sv"
  

endpackage

`endif//LVC_AHB_PKG_SV

