`ifndef RKV_AHBRAM_PKG_SV
`define RKV_AHBRAM_PKG_SV

package rkv_ahbram_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import lvc_ahb_pkg::*;
  
  `include "rkv_ahbram_reg.sv"
  `include "rkv_ahbram_config.sv"
  `include "rkv_ahbram_reg_adapter.sv"
  `include "rkv_ahbram_subscriber.sv"
  `include "rkv_ahbram_cov.sv"
  `include "rkv_ahbram_scoreboard.sv"
  `include "rkv_ahbram_virtual_sequencer.sv"
  `include "rkv_ahbram_env.sv"
  `include "rkv_ahbram_seq_lib.svh"
  `include "rkv_ahbram_tests.svh"

endpackage

`endif//RKV_AHBRAM_PKG_SV

