`ifndef RKV_AHBRAM_TESTS_SVH
`define RKV_AHBRAM_TESTS_SVH

`include "rkv_ahbram_base_test.sv"
`include "rkv_ahbram_smoke_test.sv"
`include "rkv_ahbram_diff_hsize_test.sv"
`include "rkv_ahbram_diff_haddr_test.sv"
`include "rkv_ahbram_reset_w2r_test.sv"
`include "rkv_ahbram_haddr_word_unaligned_test.sv"

`endif//RKV_AHBRAM_TESTS_SVH

