`ifndef RKV_AHBRAM_TESTS_SVH
`define RKV_AHBRAM_TESTS_SVH

`include "rkv_ahbram_base_test.sv"
`include "rkv_ahbram_smoke_test.sv"

`endif//RKV_AHBRAM_TESTS_SVH

